
// Copyright (c) 2014 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

// bsv libraries
import Vector::*;

// Connectal libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import MemTypes::*;
import MemPortal::*;
import HostInterface::*;

// generated by tool
import LedControllerRequest::*;
import SwitchRequest::*;
import SwitchIndication::*;

// defined by user
import Controller::*;
import SwitchPins::*;

module mkConnectalTop(ConnectalTop#(PhysAddrWidth,DataBusWidth,SwitchPins,0));

   // instantiate user portals
   SwitchIndicationProxy switchIndicationProxy <- mkSwitchIndicationProxy(SwitchIndicationPortal);
   Controller controller <- mkControllerRequest(switchIndicationProxy.ifc);
   
   LedControllerRequestWrapper ledControllerRequestWrapper <- mkLedControllerRequestWrapper(LedControllerRequestPortal,controller.ledRequest);
   SwitchRequestWrapper switchRequestWrapper <- mkSwitchRequestWrapper(SwitchRequestPortal,controller.switchRequest);
   
   Vector#(3,StdPortal) portals;
   portals[0] = ledControllerRequestWrapper.portalIfc;
   portals[1] = switchRequestWrapper.portalIfc;
   portals[2] = switchIndicationProxy.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = nil;
   interface pins = controller.switchPins;

endmodule : mkConnectalTop

export SwitchPins::*;
export mkConnectalTop;

